`include "params.sv"

module FloppyComp_V1 (
    input logic clock

);


    
endmodule